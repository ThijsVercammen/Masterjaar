-- Thijs Vercammen
-- r0638823
-- Digitale Synthese- labo
-- 7 segment decoder
-- November 2020
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;

entity seg_dec_r is
port (
	zevenseg_data:	in  std_logic_vector(3 downto 0);
	led:	 	out std_logic_vector(6 downto 0)
	);
end seg_dec_r;

architecture behav of seg_dec_r is
begin

comb_led_dec:PROCESS (zevenseg_data)	-- combinatorisch
BEGIN
	CASE zevenseg_data IS
    		when "0000" => led <= "0111111"; -- 0
    		when "0001" => led <= "0000110"; -- 1
    		when "0010" => led <= "1011011"; -- 2
    		when "0011" => led <= "1001111"; -- 3
    		when "0100" => led <= "1100110"; -- 4
    		when "0101" => led <= "1101101"; -- 5
    		when "0110" => led <= "1111101"; -- 6
    		when "0111" => led <= "0000111"; -- 7
    		when "1000" => led <= "1111111"; -- 8
    		when "1001" => led <= "1101111"; -- 9
    		when "1010" => led <= "1110111"; -- A
    		when "1011" => led <= "1111100"; -- b
    		when "1100" => led <= "0111001"; -- C
    		when "1101" => led <= "1011110"; -- d
    		when "1110" => led <= "1111001"; -- E
    		when "1111" => led <= "1110001"; -- F
    		when others => led <= "0000000";
	END CASE;
END PROCESS comb_led_dec;
end behav;

