-- Thijs Vercammen
-- r0638823
-- Digitale Synthese- labo
-- 7 segment decoder testbench
-- Vrijdag 24 November 2020
-- seg_dec_r_tb.vhd
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity seg_dec_r_tb is
end seg_dec_r_tb;

architecture structural of seg_dec_r_tb is 

-- Component Declaration
component seg_dec_r
port (
 	--clk: 		in std_logic;
	zevenseg_data:	in  std_logic_vector(3 downto 0):=(others => '0');
	led:	 	out std_logic_vector(6 downto 0):=(others => '0')
  );
end component;

-- uut1, uut2 verschillend initaties van component counter, handig om meerdere counters te gebruiken (ipv copy paste)
for uut : seg_dec_r use entity work.seg_dec_r(behav);
 
constant period : time := 100 ns;
constant delay  : time :=  10 ns;
signal end_of_sim : boolean := false;

-- interne testcomponent waarden, moeten niet noodzakelijk hetzelfde zijn als de entiteit
--signal clk:		std_logic;
signal zevenseg_data: std_logic_vector(3 downto 0);
signal led: std_logic_vector(6 downto 0);

BEGIN

  uut: seg_dec_r PORT MAP(
  -- links naam entiteit, rechts naam testcomponent
	--clk 		=> clk,
	zevenseg_data 	=> zevenseg_data,
	led		=> led
  );
  
tb : PROCESS
-- procedure -> functie aanmaken die kan opgeroepen worden
   procedure tbvector(constant stimvect : in std_logic_vector(3 downto 0))is
     begin
      zevenseg_data <= stimvect(3 downto 0);
      wait for period;
   end tbvector;
   BEGIN
      -- reset
      tbvector("0000");  
      tbvector("0001");
      tbvector("0010");
      tbvector("0011");
      tbvector("0100");
      tbvector("0101");
      tbvector("0110");
      tbvector("0111");
      tbvector("1000");
      tbvector("1001");
      tbvector("1010");
      tbvector("1011");
      tbvector("1100");
      tbvector("1101");
      tbvector("1110");
      tbvector("1111");
                        
      end_of_sim <= true;
      wait;
   END PROCESS;

  END;




