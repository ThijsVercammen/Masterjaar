-- Thijs Vercammen
-- r0638823
-- Digitale Synthese- labo
-- datalink testbench
-- Dinsdag 27 oktober 2020
-- datalink_tb.vhd
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity datalink_tb is
end datalink_tb;

architecture structural of datalink_tb is 

-- Component Declaration
component datalink
port (
	clk,rst:	in std_logic;
	clk_en:		in std_logic;
	pn_start:	in std_logic;
	ud_counter:	in std_logic_vector(3 downto 0):="0000";
	unencrypted:	out std_logic
  );
end component;

-- uut1, uut2 verschillend initaties van component counter, handig om meerdere counters te gebruiken (ipv copy paste)
for uut : datalink use entity work.datalink(behav);
 
constant period : time := 100 ns;
constant delay  : time :=  10 ns;
signal end_of_sim : boolean := false;

-- interne testcomponent waarden, moeten niet noodzakelijk hetzelfde zijn als de entiteit
signal clk,rst:		std_logic;
signal clk_en:		std_logic;
signal pn_start:	std_logic;
signal ud_counter:	std_logic_vector(3 downto 0):="0000";
signal unencrypted:	std_logic;

BEGIN

  uut: datalink PORT MAP(
  -- links naam entiteit, rechts naam testcomponent
	clk		=> clk,
	clk_en		=> clk_en,
	rst		=> rst,
	pn_start	=> pn_start,
	ud_counter	=> ud_counter,
	unencrypted	=> unencrypted
  );

  clock : process
   begin 
       clk <= '0';
       wait for period/2;
     loop
       clk <= '0';
       wait for period/2;
       clk <= '1';
       wait for period/2;
       exit when end_of_sim;
     end loop;
     wait;
   end process clock;
  
tb : PROCESS
-- procedure -> functie aanmaken die kan opgeroepen worden
   procedure tbvector(constant stimvect : in std_logic_vector(5 downto 0))is
     begin
      ud_counter <= stimvect(5 downto 2);
      pn_start <= stimvect(1);
      rst <= stimvect(0);
      clk_en <= '1';
      wait for period;
   end tbvector;
   BEGIN
      -- reset
      tbvector("000001");
      tbvector("000001");
      
      -- counting
      tbvector("101010"); -- up 1
      wait for period*15;
      
      tbvector("001110"); -- up 3
      wait for period*15;

      tbvector("110010"); -- up 3
      wait for period*5;

      tbvector("110110"); -- up 3
      wait for period*20;

      tbvector("000001"); -- reset
      tbvector("000001"); -- reset
                       
      end_of_sim <= true;
      wait;
   END PROCESS;

  END;
